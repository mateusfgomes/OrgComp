LIBRARY IEEE;
USE  IEEE.STD_LOGIC_1164.ALL;
USE  IEEE.STD_LOGIC_ARITH.ALL;
USE  IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY hex_2_7seg IS
	PORT(
			HEX : IN STD_LOGIC_VECTOR(3 downto 0);
			SEG : OUT STD_LOGIC_VECTOR(6 DOWNTO 0)
		);
END hex_2_7seg;

ARCHITECTURE main OF hex_2_7seg IS
SIGNAL SEG_DATA : STD_LOGIC_VECTOR(6 DOWNTO 0);
BEGIN
	PROCESS(HEX)
	BEGIN
		CASE HEX IS
			WHEN "0000" =>
				SEG_DATA <= "0111111";
			WHEN "0001" =>
				SEG_DATA <= "0000110";
			WHEN "0010" =>
				SEG_DATA <= "1011011";
			WHEN "0011" =>
				SEG_DATA <= "1001111";
			WHEN "0100" =>
				SEG_DATA <= "1100110";
			WHEN "0101" =>
				SEG_DATA <= "1101101";
			WHEN "0110" =>
				SEG_DATA <= "1111101";
			WHEN "0111" =>
				SEG_DATA <= "0000111";
			WHEN "1000" =>
				SEG_DATA <= "1111111";
			WHEN "1001" =>
				SEG_DATA <= "1101111"; 
			WHEN "1010" =>
				SEG_DATA <= "1110111";
			WHEN "1011" =>
				SEG_DATA <= "1111100"; 
			WHEN "1100" =>
				SEG_DATA <= "0111001"; 
			WHEN "1101" =>
				SEG_DATA <= "1011110"; 
			WHEN "1110" =>
				SEG_DATA <= "1111001"; 
			WHEN "1111" =>
				SEG_DATA <= "1110001"; 
			WHEN OTHERS =>
				SEG_DATA <= "1000000";
		END CASE;
	END PROCESS;

SEG <= NOT SEG_DATA;

END main;