LIBRARY IEEE;
USE  IEEE.STD_LOGIC_1164.all;
USE  IEEE.STD_LOGIC_ARITH.all;
USE  IEEE.STD_LOGIC_UNSIGNED.all;

ENTITY KB_RECEIVER IS
	PORT(	CLK		: IN STD_LOGIC;
			RST		: IN STD_LOGIC;
			KBCLK		: IN STD_LOGIC;
			KBDATA	: IN STD_LOGIC;
			
			KEYSTATE : OUT STD_LOGIC;
			KEY		: OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
			EXTENDED : OUT STD_LOGIC
		);
END KB_RECEIVER;

ARCHITECTURE main OF KB_RECEIVER IS

	SIGNAL KBCLKF : STD_LOGIC;

BEGIN
	PROCESS(KBCLKF, RST)
	
		VARIABLE REC_DATA 	: STD_LOGIC_VECTOR(7 DOWNTO 0);
		VARIABLE STATE 		: STD_LOGIC_VECTOR(3 DOWNTO 0);
		VARIABLE ITERATOR 	: INTEGER RANGE 0 TO 10;
		VARIABLE UNPRESSING	: STD_LOGIC;
		
	BEGIN
		IF(RST = '1') THEN
			STATE 		:= x"0";
			ITERATOR 	:= 0;
			UNPRESSING 	:= '0';
			KEY 			<= x"FF";
			KEYSTATE 	<= '0';
			EXTENDED 	<= '0';
		ELSIF(KBCLKF'EVENT AND KBCLKF = '0') THEN
		
			CASE STATE IS
			
				WHEN x"0" =>
					KEYSTATE <= '1';
					STATE := x"1";
					
				-- carrega rec_data com 8 bits vindos do teclado
				-- cada bit chega em um pulso do clock
				WHEN x"1" =>
					REC_DATA(ITERATOR)	:= KBDATA;
					ITERATOR					:= ITERATOR + 1;
					IF(ITERATOR = 8) THEN
						STATE := x"2";
					END IF;
					
				WHEN x"2" =>
					IF(REC_DATA = x"E0") THEN
						EXTENDED <= '1';
					ELSIF(REC_DATA = x"F0") THEN
						UNPRESSING := '1';
					ELSIF(UNPRESSING = '1') THEN
						UNPRESSING := '0';
						KEYSTATE <= '0';
						EXTENDED <= '0';
						KEY <= x"FF";
					ELSE
						KEY <= REC_DATA;
					END IF;
					ITERATOR := 0;
					STATE := x"3";
					
				WHEN x"3" =>
					STATE := x"0";
					
				WHEN OTHERS =>
				
			END CASE;
		END IF;
	END PROCESS;

	PROCESS(CLK)
	
		VARIABLE CLK_FILTER : STD_LOGIC_VECTOR(7 DOWNTO 0);
		
	BEGIN
		IF(CLK'EVENT AND CLK = '1') THEN
			CLK_FILTER(6 DOWNTO 0) := CLK_FILTER(7 DOWNTO 1); -- shifta para a direita
			CLK_FILTER(7) := KBCLK;
			IF(CLK_FILTER = "11111111") THEN
				KBCLKF <= '1';
			ELSIF(CLK_FILTER = "00000000") THEN 
				KBCLKF <= '0';
			END IF;
		END IF;
	END PROCESS;
END main;